magic
tech sky130A
magscale 1 2
timestamp 1671535159
<< nwell >>
rect 1066 116677 178886 117243
rect 1066 115589 178886 116155
rect 1066 114501 178886 115067
rect 1066 113413 178886 113979
rect 1066 112325 178886 112891
rect 1066 111237 178886 111803
rect 1066 110149 178886 110715
rect 1066 109061 178886 109627
rect 1066 107973 178886 108539
rect 1066 106885 178886 107451
rect 1066 105797 178886 106363
rect 1066 104709 178886 105275
rect 1066 103621 178886 104187
rect 1066 102533 178886 103099
rect 1066 101445 178886 102011
rect 1066 100357 178886 100923
rect 1066 99269 178886 99835
rect 1066 98181 178886 98747
rect 1066 97093 178886 97659
rect 1066 96005 178886 96571
rect 1066 94917 178886 95483
rect 1066 93829 178886 94395
rect 1066 92741 178886 93307
rect 1066 91653 178886 92219
rect 1066 90565 178886 91131
rect 1066 89477 178886 90043
rect 1066 88389 178886 88955
rect 1066 87301 178886 87867
rect 1066 86213 178886 86779
rect 1066 85125 178886 85691
rect 1066 84037 178886 84603
rect 1066 82949 178886 83515
rect 1066 81861 178886 82427
rect 1066 80773 178886 81339
rect 1066 79685 178886 80251
rect 1066 78597 178886 79163
rect 1066 77509 178886 78075
rect 1066 76421 178886 76987
rect 1066 75333 178886 75899
rect 1066 74245 178886 74811
rect 1066 73157 178886 73723
rect 1066 72069 178886 72635
rect 1066 70981 178886 71547
rect 1066 69893 178886 70459
rect 1066 68805 178886 69371
rect 1066 67717 178886 68283
rect 1066 66629 178886 67195
rect 1066 65541 178886 66107
rect 1066 64453 178886 65019
rect 1066 63365 178886 63931
rect 1066 62277 178886 62843
rect 1066 61189 178886 61755
rect 1066 60101 178886 60667
rect 1066 59013 178886 59579
rect 1066 57925 178886 58491
rect 1066 56837 178886 57403
rect 1066 55749 178886 56315
rect 1066 54661 178886 55227
rect 1066 53573 178886 54139
rect 1066 52485 178886 53051
rect 1066 51397 178886 51963
rect 1066 50309 178886 50875
rect 1066 49221 178886 49787
rect 1066 48133 178886 48699
rect 1066 47045 178886 47611
rect 1066 45957 178886 46523
rect 1066 44869 178886 45435
rect 1066 43781 178886 44347
rect 1066 42693 178886 43259
rect 1066 41605 178886 42171
rect 1066 40517 178886 41083
rect 1066 39429 178886 39995
rect 1066 38341 178886 38907
rect 1066 37253 178886 37819
rect 1066 36165 178886 36731
rect 1066 35077 178886 35643
rect 1066 33989 178886 34555
rect 1066 32901 178886 33467
rect 1066 31813 178886 32379
rect 1066 30725 178886 31291
rect 1066 29637 178886 30203
rect 1066 28549 178886 29115
rect 1066 27461 178886 28027
rect 1066 26373 178886 26939
rect 1066 25285 178886 25851
rect 1066 24197 178886 24763
rect 1066 23109 178886 23675
rect 1066 22021 178886 22587
rect 1066 20933 178886 21499
rect 1066 19845 178886 20411
rect 1066 18757 178886 19323
rect 1066 17669 178886 18235
rect 1066 16581 178886 17147
rect 1066 15493 178886 16059
rect 1066 14405 178886 14971
rect 1066 13317 178886 13883
rect 1066 12229 178886 12795
rect 1066 11141 178886 11707
rect 1066 10053 178886 10619
rect 1066 8965 178886 9531
rect 1066 7877 178886 8443
rect 1066 6789 178886 7355
rect 1066 5701 178886 6267
rect 1066 4613 178886 5179
rect 1066 3525 178886 4091
rect 1066 2437 178886 3003
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 1104 1708 178848 117552
<< metal2 >>
rect 2042 0 2098 800
rect 5630 0 5686 800
rect 9218 0 9274 800
rect 12806 0 12862 800
rect 16394 0 16450 800
rect 19982 0 20038 800
rect 23570 0 23626 800
rect 27158 0 27214 800
rect 30746 0 30802 800
rect 34334 0 34390 800
rect 37922 0 37978 800
rect 41510 0 41566 800
rect 45098 0 45154 800
rect 48686 0 48742 800
rect 52274 0 52330 800
rect 55862 0 55918 800
rect 59450 0 59506 800
rect 63038 0 63094 800
rect 66626 0 66682 800
rect 70214 0 70270 800
rect 73802 0 73858 800
rect 77390 0 77446 800
rect 80978 0 81034 800
rect 84566 0 84622 800
rect 88154 0 88210 800
rect 91742 0 91798 800
rect 95330 0 95386 800
rect 98918 0 98974 800
rect 102506 0 102562 800
rect 106094 0 106150 800
rect 109682 0 109738 800
rect 113270 0 113326 800
rect 116858 0 116914 800
rect 120446 0 120502 800
rect 124034 0 124090 800
rect 127622 0 127678 800
rect 131210 0 131266 800
rect 134798 0 134854 800
rect 138386 0 138442 800
rect 141974 0 142030 800
rect 145562 0 145618 800
rect 149150 0 149206 800
rect 152738 0 152794 800
rect 156326 0 156382 800
rect 159914 0 159970 800
rect 163502 0 163558 800
rect 167090 0 167146 800
rect 170678 0 170734 800
rect 174266 0 174322 800
rect 177854 0 177910 800
<< obsm2 >>
rect 2044 856 177908 117541
rect 2154 734 5574 856
rect 5742 734 9162 856
rect 9330 734 12750 856
rect 12918 734 16338 856
rect 16506 734 19926 856
rect 20094 734 23514 856
rect 23682 734 27102 856
rect 27270 734 30690 856
rect 30858 734 34278 856
rect 34446 734 37866 856
rect 38034 734 41454 856
rect 41622 734 45042 856
rect 45210 734 48630 856
rect 48798 734 52218 856
rect 52386 734 55806 856
rect 55974 734 59394 856
rect 59562 734 62982 856
rect 63150 734 66570 856
rect 66738 734 70158 856
rect 70326 734 73746 856
rect 73914 734 77334 856
rect 77502 734 80922 856
rect 81090 734 84510 856
rect 84678 734 88098 856
rect 88266 734 91686 856
rect 91854 734 95274 856
rect 95442 734 98862 856
rect 99030 734 102450 856
rect 102618 734 106038 856
rect 106206 734 109626 856
rect 109794 734 113214 856
rect 113382 734 116802 856
rect 116970 734 120390 856
rect 120558 734 123978 856
rect 124146 734 127566 856
rect 127734 734 131154 856
rect 131322 734 134742 856
rect 134910 734 138330 856
rect 138498 734 141918 856
rect 142086 734 145506 856
rect 145674 734 149094 856
rect 149262 734 152682 856
rect 152850 734 156270 856
rect 156438 734 159858 856
rect 160026 734 163446 856
rect 163614 734 167034 856
rect 167202 734 170622 856
rect 170790 734 174210 856
rect 174378 734 177798 856
<< obsm3 >>
rect 4210 1939 173486 117537
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 15515 2211 19488 40085
rect 19968 2211 34848 40085
rect 35328 2211 50208 40085
rect 50688 2211 65568 40085
rect 66048 2211 80928 40085
rect 81408 2211 82005 40085
<< labels >>
rlabel metal2 s 9218 0 9274 800 6 clk
port 1 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 execute
port 2 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 input_val[0]
port 3 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 input_val[1]
port 4 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 input_val[2]
port 5 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 input_val[3]
port 6 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 input_val[4]
port 7 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 input_val[5]
port 8 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 input_val[6]
port 9 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 input_val[7]
port 10 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 io_oeb[0]
port 11 nsew signal output
rlabel metal2 s 156326 0 156382 800 6 io_oeb[10]
port 12 nsew signal output
rlabel metal2 s 159914 0 159970 800 6 io_oeb[11]
port 13 nsew signal output
rlabel metal2 s 163502 0 163558 800 6 io_oeb[12]
port 14 nsew signal output
rlabel metal2 s 167090 0 167146 800 6 io_oeb[13]
port 15 nsew signal output
rlabel metal2 s 170678 0 170734 800 6 io_oeb[14]
port 16 nsew signal output
rlabel metal2 s 174266 0 174322 800 6 io_oeb[15]
port 17 nsew signal output
rlabel metal2 s 177854 0 177910 800 6 io_oeb[16]
port 18 nsew signal output
rlabel metal2 s 124034 0 124090 800 6 io_oeb[1]
port 19 nsew signal output
rlabel metal2 s 127622 0 127678 800 6 io_oeb[2]
port 20 nsew signal output
rlabel metal2 s 131210 0 131266 800 6 io_oeb[3]
port 21 nsew signal output
rlabel metal2 s 134798 0 134854 800 6 io_oeb[4]
port 22 nsew signal output
rlabel metal2 s 138386 0 138442 800 6 io_oeb[5]
port 23 nsew signal output
rlabel metal2 s 141974 0 142030 800 6 io_oeb[6]
port 24 nsew signal output
rlabel metal2 s 145562 0 145618 800 6 io_oeb[7]
port 25 nsew signal output
rlabel metal2 s 149150 0 149206 800 6 io_oeb[8]
port 26 nsew signal output
rlabel metal2 s 152738 0 152794 800 6 io_oeb[9]
port 27 nsew signal output
rlabel metal2 s 2042 0 2098 800 6 reset
port 28 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 result[0]
port 29 nsew signal output
rlabel metal2 s 95330 0 95386 800 6 result[10]
port 30 nsew signal output
rlabel metal2 s 98918 0 98974 800 6 result[11]
port 31 nsew signal output
rlabel metal2 s 102506 0 102562 800 6 result[12]
port 32 nsew signal output
rlabel metal2 s 106094 0 106150 800 6 result[13]
port 33 nsew signal output
rlabel metal2 s 109682 0 109738 800 6 result[14]
port 34 nsew signal output
rlabel metal2 s 113270 0 113326 800 6 result[15]
port 35 nsew signal output
rlabel metal2 s 116858 0 116914 800 6 result[16]
port 36 nsew signal output
rlabel metal2 s 63038 0 63094 800 6 result[1]
port 37 nsew signal output
rlabel metal2 s 66626 0 66682 800 6 result[2]
port 38 nsew signal output
rlabel metal2 s 70214 0 70270 800 6 result[3]
port 39 nsew signal output
rlabel metal2 s 73802 0 73858 800 6 result[4]
port 40 nsew signal output
rlabel metal2 s 77390 0 77446 800 6 result[5]
port 41 nsew signal output
rlabel metal2 s 80978 0 81034 800 6 result[6]
port 42 nsew signal output
rlabel metal2 s 84566 0 84622 800 6 result[7]
port 43 nsew signal output
rlabel metal2 s 88154 0 88210 800 6 result[8]
port 44 nsew signal output
rlabel metal2 s 91742 0 91798 800 6 result[9]
port 45 nsew signal output
rlabel metal2 s 12806 0 12862 800 6 sel_in[0]
port 46 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 sel_in[1]
port 47 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 sel_in[2]
port 48 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 sel_out[0]
port 49 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 sel_out[1]
port 50 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 51 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 51 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 51 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 51 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 51 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 51 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 52 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 52 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 52 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 52 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 52 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 16686316
string GDS_FILE /home/radhe/opensource/matrix_multiply_mpw8/openlane/matrix_multiply/runs/22_12_20_16_32/results/signoff/matrix_multiply.magic.gds
string GDS_START 886320
<< end >>

